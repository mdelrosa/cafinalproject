//master module to handle switching between modes

module master(
	input switch
	input clk
	output mode
);